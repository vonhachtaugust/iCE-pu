-------------------------------------------------------------------------------
-- Title      : icePU package
-- Project    : icePU
-------------------------------------------------------------------------------
-- File       : icePU_pkg.vhdl
-- Author     : August  <vonhachtaugust@gmail.com>
-- Company    :
-- Created    : 2020-07-01
-- Last update: 2020-07-07
-- Platform   : Lattice iCEstick Evaluation Kit
-- Standard   : VHDL'08
-------------------------------------------------------------------------------
-- Description: icePU package
-------------------------------------------------------------------------------
-- Copyright (c) 2020
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2020-07-01  1.0      August  Created
-------------------------------------------------------------------------------

package icePU_pkg is

  -- Constants
  -- Types
  -- Functions

end package icePU_pkg;

package body icePU_pkg is

  -- Functions

end package body icePu_pkg;