-------------------------------------------------------------------------------
-- Title      : Register file test bench
-- Project    : icePU
-------------------------------------------------------------------------------
-- File       : reg32_8_tb.vhdl
-- Author     : August  <vonhachtaugust@gmail.com>
-- Company    :
-- Created    : 2020-07-01
-- Last update: 2020-07-07
-- Platform   : Lattice iCEstick Evaluation Kit
-- Standard   : VHDL'08
-------------------------------------------------------------------------------
-- Description: Register file test bench
-------------------------------------------------------------------------------
-- Copyright (c) 2020
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2020-07-01  1.0      August  Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity reg32_8_tb is
end entity reg32_8_tb;

architecture rtl of reg32_8 is
begin
end architecture rtl;